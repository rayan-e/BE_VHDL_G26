COMPONENT traitement 
	port(
		clk : in std_logic;
		cs_in : in std_logic;
		Cs :out std_logic;
		debut_coverstion : in std_logic;
		reset : in std_logic;
		data_in : in std_logic;
		data_out : out std_logic_vector(11 downto 0)
		);
END COMPONENT;